	mem(0) := To_stdlogicvector(X"01");
	mem(1) := To_stdlogicvector(X"F0");
	mem(2) := To_stdlogicvector(X"04");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"03");
	mem(5) := To_stdlogicvector(X"15");
	mem(6) := To_stdlogicvector(X"C0");
	mem(7) := To_stdlogicvector(X"C1");
	mem(8) := To_stdlogicvector(X"10");
	mem(9) := To_stdlogicvector(X"2C");
	mem(10) := To_stdlogicvector(X"11");
	mem(11) := To_stdlogicvector(X"2E");
	mem(12) := To_stdlogicvector(X"12");
	mem(13) := To_stdlogicvector(X"3C");
	mem(14) := To_stdlogicvector(X"13");
	mem(15) := To_stdlogicvector(X"3E");
	mem(16) := To_stdlogicvector(X"0D");
	mem(17) := To_stdlogicvector(X"60");
	mem(20) := To_stdlogicvector(X"0D");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"60");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"A5");
	mem(25) := To_stdlogicvector(X"13");
	mem(26) := To_stdlogicvector(X"65");
	mem(27) := To_stdlogicvector(X"12");
	mem(28) := To_stdlogicvector(X"7D");
	mem(29) := To_stdlogicvector(X"12");
	mem(30) := To_stdlogicvector(X"65");
	mem(31) := To_stdlogicvector(X"52");
	mem(32) := To_stdlogicvector(X"63");
	mem(33) := To_stdlogicvector(X"D4");
	mem(34) := To_stdlogicvector(X"93");
	mem(35) := To_stdlogicvector(X"D4");
	mem(36) := To_stdlogicvector(X"21");
	mem(37) := To_stdlogicvector(X"F0");
	mem(38) := To_stdlogicvector(X"B4");
	mem(39) := To_stdlogicvector(X"D4");
	mem(40) := To_stdlogicvector(X"0C");
	mem(41) := To_stdlogicvector(X"E0");
	mem(42) := To_stdlogicvector(X"0E");
	mem(43) := To_stdlogicvector(X"48");
	mem(44) := To_stdlogicvector(X"00");
	mem(45) := To_stdlogicvector(X"C0");
	mem(46) := To_stdlogicvector(X"16");
	mem(47) := To_stdlogicvector(X"04");
	mem(48) := To_stdlogicvector(X"C0");
	mem(49) := To_stdlogicvector(X"C1");
	mem(50) := To_stdlogicvector(X"06");
	mem(51) := To_stdlogicvector(X"12");
	mem(52) := To_stdlogicvector(X"7F");
	mem(53) := To_stdlogicvector(X"9B");
	mem(54) := To_stdlogicvector(X"45");
	mem(55) := To_stdlogicvector(X"12");
	mem(56) := To_stdlogicvector(X"46");
	mem(57) := To_stdlogicvector(X"16");
	mem(58) := To_stdlogicvector(X"00");
	mem(59) := To_stdlogicvector(X"00");
	mem(60) := To_stdlogicvector(X"01");
	mem(61) := To_stdlogicvector(X"00");
	mem(62) := To_stdlogicvector(X"05");
	mem(63) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"01");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"80");
	mem(67) := To_stdlogicvector(X"14");
	mem(68) := To_stdlogicvector(X"45");
	mem(69) := To_stdlogicvector(X"12");
	mem(70) := To_stdlogicvector(X"FD");
	mem(71) := To_stdlogicvector(X"0B");
	mem(72) := To_stdlogicvector(X"86");
	mem(73) := To_stdlogicvector(X"1E");
	mem(74) := To_stdlogicvector(X"86");
	mem(75) := To_stdlogicvector(X"54");
	mem(76) := To_stdlogicvector(X"C5");
	mem(77) := To_stdlogicvector(X"16");
	mem(78) := To_stdlogicvector(X"07");
	mem(79) := To_stdlogicvector(X"04");
	mem(80) := To_stdlogicvector(X"C6");
	mem(81) := To_stdlogicvector(X"12");
	mem(82) := To_stdlogicvector(X"C6");
	mem(83) := To_stdlogicvector(X"11");
	mem(84) := To_stdlogicvector(X"02");
	mem(85) := To_stdlogicvector(X"14");
	mem(86) := To_stdlogicvector(X"45");
	mem(87) := To_stdlogicvector(X"12");
	mem(88) := To_stdlogicvector(X"FD");
	mem(89) := To_stdlogicvector(X"0B");
	mem(90) := To_stdlogicvector(X"F6");
	mem(91) := To_stdlogicvector(X"0F");
	mem(92) := To_stdlogicvector(X"9E");
	mem(93) := To_stdlogicvector(X"6F");
	mem(94) := To_stdlogicvector(X"FF");
	mem(95) := To_stdlogicvector(X"0F");
