--
-- VHDL Architecture ece411.mp3_IR.untitled
--
-- Created:
--          by - hwoods2.ece411_G3 (gllnx11.ews.illinois.edu)
--          at - 17:32:36 10/20/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY mp3_IR IS
   PORT(
      LoadIR      : IN     std_logic;
      instruction : IN     LC3b_word;
      clk         : IN     std_logic;
      Opcode      : OUT    LC3b_opcode;
      SrcA        : OUT    LC3b_reg;
      SrcB        : OUT    LC3b_reg;
      destin      : OUT    LC3b_reg;
      index6      : OUT    LC3b_index6;
      offset9     : OUT    LC3b_offset9;
      reset_l     : IN     std_logic
   );

-- Declarations

END mp3_IR ;

--
ARCHITECTURE untitled OF mp3_IR IS
BEGIN
  ------------------------------
  VHDL_REG_IR : PROCESS (CLK, LOADIR, instruction)
  ------------------------------
  BEGIN
	  IF (CLK'EVENT AND (CLK = '1') AND (CLK'LAST_VALUE = '0')) THEN
		  IF (LOADIR = '1') THEN
			  VAL_IR <= MDROUT AFTER DELAY_REG;
		  END IF;
	  END IF;
  END PROCESS VHDL_REG_IR;
  OPCODE <= VAL_IR(15 DOWNTO 12);
  SRCA <= VAL_IR(8 DOWNTO 6);
  SRCB <= VAL_IR(2 DOWNTO 0);
  Destin <= VAL_IR(11 DOWNTO 9);
  OFFSET9 <= VAL_IR(8 DOWNTO 0);
  INDEX6 <= VAL_IR(5 DOWNTO 0);
  
END ARCHITECTURE untitled;

