--
-- VHDL Architecture ece411.mp3_Control.untitled
--
-- Created:
--          by - hwoods2.ece411_G3 (gllnx11.ews.illinois.edu)
--          at - 17:17:12 10/20/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY mp3_Control IS
   PORT( 
      clk : IN     std_logic
   );

-- Declarations

END mp3_Control ;

--
ARCHITECTURE untitled OF mp3_Control IS
BEGIN
END ARCHITECTURE untitled;

