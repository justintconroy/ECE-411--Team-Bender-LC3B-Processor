	mem(0) := To_stdlogicvector(X"25");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"25");
	mem(3) := To_stdlogicvector(X"14");
	mem(4) := To_stdlogicvector(X"81");
	mem(5) := To_stdlogicvector(X"12");
	mem(6) := To_stdlogicvector(X"BF");
	mem(7) := To_stdlogicvector(X"14");
	mem(8) := To_stdlogicvector(X"09");
	mem(9) := To_stdlogicvector(X"74");
	mem(10) := To_stdlogicvector(X"05");
	mem(11) := To_stdlogicvector(X"48");
	mem(12) := To_stdlogicvector(X"09");
	mem(13) := To_stdlogicvector(X"E8");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"41");
	mem(16) := To_stdlogicvector(X"FF");
	mem(17) := To_stdlogicvector(X"0F");
	mem(18) := To_stdlogicvector(X"DD");
	mem(19) := To_stdlogicvector(X"DD");
	mem(20) := To_stdlogicvector(X"FF");
	mem(21) := To_stdlogicvector(X"FF");
	mem(22) := To_stdlogicvector(X"0A");
	mem(23) := To_stdlogicvector(X"6A");
	mem(24) := To_stdlogicvector(X"64");
	mem(25) := To_stdlogicvector(X"DB");
	mem(26) := To_stdlogicvector(X"74");
	mem(27) := To_stdlogicvector(X"DB");
	mem(28) := To_stdlogicvector(X"54");
	mem(29) := To_stdlogicvector(X"DB");
	mem(30) := To_stdlogicvector(X"C0");
	mem(31) := To_stdlogicvector(X"C1");
	mem(32) := To_stdlogicvector(X"0A");
	mem(33) := To_stdlogicvector(X"62");
	mem(34) := To_stdlogicvector(X"61");
	mem(35) := To_stdlogicvector(X"12");
	mem(36) := To_stdlogicvector(X"81");
	mem(37) := To_stdlogicvector(X"12");
	mem(38) := To_stdlogicvector(X"42");
	mem(39) := To_stdlogicvector(X"52");
	mem(40) := To_stdlogicvector(X"61");
	mem(41) := To_stdlogicvector(X"D2");
	mem(42) := To_stdlogicvector(X"F2");
	mem(43) := To_stdlogicvector(X"E3");
	mem(44) := To_stdlogicvector(X"09");
	mem(45) := To_stdlogicvector(X"6C");
	mem(46) := To_stdlogicvector(X"40");
	mem(47) := To_stdlogicvector(X"C0");
