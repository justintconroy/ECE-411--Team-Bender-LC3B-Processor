--
-- VHDL Architecture ece411.RipRFABit0.untitled
--
-- Created:
--          by - hwoods2.stdt (eelnx35.ews.illinois.edu)
--          at - 19:54:34 09/16/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY RipRFABit0 IS
   PORT( 
      ALUout       : IN     LC3b_word;
      clk           : IN     std_logic;
      RipRFABit0out : OUT    std_logic
   );

-- Declarations

END RipRFABit0 ;

--
ARCHITECTURE untitled OF RipRFABit0 IS
BEGIN
  RipRFABit0out <= ALUout(0);
END ARCHITECTURE untitled;

