	MEM(0) := TO_STDLOGICVECTOR(X"11");
		MEM(1) := TO_STDLOGICVECTOR(X"62");
		MEM(2) := TO_STDLOGICVECTOR(X"12");
		MEM(3) := TO_STDLOGICVECTOR(X"64");
		MEM(4) := TO_STDLOGICVECTOR(X"13");
		MEM(5) := TO_STDLOGICVECTOR(X"66");
		MEM(6) := TO_STDLOGICVECTOR(X"C2");
		MEM(7) := TO_STDLOGICVECTOR(X"18");
		MEM(8) := TO_STDLOGICVECTOR(X"C3");
		MEM(9) := TO_STDLOGICVECTOR(X"16");
		MEM(10) := TO_STDLOGICVECTOR(X"BF");
		MEM(11) := TO_STDLOGICVECTOR(X"9A");
		MEM(12) := TO_STDLOGICVECTOR(X"41");
		MEM(13) := TO_STDLOGICVECTOR(X"1B");
		MEM(14) := TO_STDLOGICVECTOR(X"05");
		MEM(15) := TO_STDLOGICVECTOR(X"19");
		MEM(16) := TO_STDLOGICVECTOR(X"FB");
		MEM(17) := TO_STDLOGICVECTOR(X"07");
		MEM(18) := TO_STDLOGICVECTOR(X"C4");
		MEM(19) := TO_STDLOGICVECTOR(X"5E");
		MEM(20) := TO_STDLOGICVECTOR(X"14");
		MEM(21) := TO_STDLOGICVECTOR(X"7E");
		MEM(22) := TO_STDLOGICVECTOR(X"14");
		MEM(23) := TO_STDLOGICVECTOR(X"62");
		MEM(24) := TO_STDLOGICVECTOR(X"FF");
		MEM(25) := TO_STDLOGICVECTOR(X"91");
		MEM(26) := TO_STDLOGICVECTOR(X"40");
		MEM(27) := TO_STDLOGICVECTOR(X"50");
		MEM(28) := TO_STDLOGICVECTOR(X"14");
		MEM(29) := TO_STDLOGICVECTOR(X"70");
		MEM(30) := TO_STDLOGICVECTOR(X"15");
		MEM(31) := TO_STDLOGICVECTOR(X"62");
		MEM(32) := TO_STDLOGICVECTOR(X"FF");
		MEM(33) := TO_STDLOGICVECTOR(X"0F");
		MEM(34) := TO_STDLOGICVECTOR(X"01");
		MEM(35) := TO_STDLOGICVECTOR(X"00");
		MEM(36) := TO_STDLOGICVECTOR(X"02");
		MEM(37) := TO_STDLOGICVECTOR(X"00");
		MEM(38) := TO_STDLOGICVECTOR(X"08");
		MEM(39) := TO_STDLOGICVECTOR(X"00");
		MEM(40) := TO_STDLOGICVECTOR(X"00");
		MEM(41) := TO_STDLOGICVECTOR(X"00");
		MEM(42) := TO_STDLOGICVECTOR(X"0D");
		MEM(43) := TO_STDLOGICVECTOR(X"60");
