	mem(0) := To_stdlogicvector(X"97");
	mem(1) := To_stdlogicvector(X"61");
	mem(2) := To_stdlogicvector(X"11");
	mem(3) := To_stdlogicvector(X"04");
	mem(4) := To_stdlogicvector(X"06");
	mem(5) := To_stdlogicvector(X"12");
	mem(6) := To_stdlogicvector(X"7F");
	mem(7) := To_stdlogicvector(X"9B");
	mem(8) := To_stdlogicvector(X"45");
	mem(9) := To_stdlogicvector(X"12");
	mem(10) := To_stdlogicvector(X"46");
	mem(11) := To_stdlogicvector(X"16");
	mem(12) := To_stdlogicvector(X"80");
	mem(13) := To_stdlogicvector(X"14");
	mem(14) := To_stdlogicvector(X"45");
	mem(15) := To_stdlogicvector(X"12");
	mem(16) := To_stdlogicvector(X"FD");
	mem(17) := To_stdlogicvector(X"0B");
	mem(18) := To_stdlogicvector(X"86");
	mem(19) := To_stdlogicvector(X"1E");
	mem(20) := To_stdlogicvector(X"86");
	mem(21) := To_stdlogicvector(X"54");
	mem(22) := To_stdlogicvector(X"C5");
	mem(23) := To_stdlogicvector(X"16");
	mem(24) := To_stdlogicvector(X"07");
	mem(25) := To_stdlogicvector(X"04");
	mem(26) := To_stdlogicvector(X"C6");
	mem(27) := To_stdlogicvector(X"12");
	mem(28) := To_stdlogicvector(X"C6");
	mem(29) := To_stdlogicvector(X"11");
	mem(30) := To_stdlogicvector(X"02");
	mem(31) := To_stdlogicvector(X"14");
	mem(32) := To_stdlogicvector(X"45");
	mem(33) := To_stdlogicvector(X"12");
	mem(34) := To_stdlogicvector(X"FD");
	mem(35) := To_stdlogicvector(X"0B");
	mem(36) := To_stdlogicvector(X"F6");
	mem(37) := To_stdlogicvector(X"0F");
	mem(38) := To_stdlogicvector(X"96");
	mem(39) := To_stdlogicvector(X"6F");
	mem(40) := To_stdlogicvector(X"FF");
	mem(41) := To_stdlogicvector(X"0F");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"01");
	mem(45) := To_stdlogicvector(X"00");
	mem(46) := To_stdlogicvector(X"05");
	mem(47) := To_stdlogicvector(X"00");
