--
-- VHDL Architecture ece411.dirtydelay.untitled
--
-- Created:
--          by - hwoods2.stdt (gllnx26.ews.illinois.edu)
--          at - 00:27:55 10/08/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY dirtydelay IS
-- Declarations

END dirtydelay ;

--
ARCHITECTURE untitled OF dirtydelay IS
BEGIN
END ARCHITECTURE untitled;

