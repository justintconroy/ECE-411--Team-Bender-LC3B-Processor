--
-- VHDL Architecture ece411.BRadd.untitled
--
-- Created:
--          by - hwoods2.stdt (eelnx29.ews.illinois.edu)
--          at - 16:22:09 08/30/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY BRadd IS
   PORT( 
      ADJ9out  : IN     LC3b_word;
      PCout    : IN     LC3b_word;
      clk      : IN     std_logic;
      BRaddout : OUT    LC3b_word
   );

-- Declarations

END BRadd ;

--
ARCHITECTURE untitled OF BRadd IS
BEGIN
  VHDL_BRadd : PROCESS (ADJ9out, PCOUT)
  BEGIN  -- PROCESS
   BRaddout <= STD_LOGIC_VECTOR(UNSIGNED(PCOUT) + UNSIGNED(ADJ9out)) AFTER DELAY_ADDER;
  END PROCESS;
END ARCHITECTURE untitled;

