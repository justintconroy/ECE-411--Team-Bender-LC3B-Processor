--
-- VHDL Architecture ece411.Way.untitled
--
-- Created:
--          by - hwoods2.stdt (eelnx28.ews.illinois.edu)
--          at - 16:06:03 09/25/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Way IS
   PORT( 
      RESET_L   : IN     std_logic;
      DataWrite : IN     std_logic;
      Index     : IN     LC3b_index;
      DataIn    : IN     LC3b_oword;
      TagIN     : IN     LC3b_tag;
      DirtyIn   : IN     std_logic;
      DataOut   : OUT    LC3b_oword;
      TagOut    : OUT    LC3b_tag;
      DirtyOut  : OUT    std_logic;
      ValidOut  : OUT    std_logic
   );

-- Declarations

END Way ;

--
ARCHITECTURE untitled OF Way IS
  	TYPE DataArray IS	array (7 downto 0) of LC3b_oword;
  	TYPE ValidArray IS array (7 downto 0) of std_logic;
  	TYPE DirtyArray IS array (7 downto 0) of std_logic;
  	TYPE TagArray IS array (7 downto 0) of LC3b_tag;
	 SIGNAL Data  : DataArray;
	 SIGNAL Valid : ValidArray;
	 SIGNAl Tag   : TagArray;
	 SIGNAL Dirty : DirtyArray;
  
   BEGIN
     --------------------------------------------------------------
		     ReadFromDataArray : PROCESS (Data, Index, Tag, Dirty, Valid)
		     --------------------------------------------------------------
         
			     VARIABLE DataIndex : integer;
			     BEGIN
				     DataIndex := to_integer(unsigned(Index));
				     DataOut  <= Data(DataIndex)  after 20 ns;
				     TagOut   <= Tag(DataIndex)   after 20 ns;
				     DirtyOut <= Dirty(DataIndex) after 20 ns;
				     ValidOut <= Valid(DataIndex) after 20 ns;
		         
		     END PROCESS ReadFromDataArray;
	     
		     --------------------------------------------------------------
		     WriteToDataArray : PROCESS (RESET_L, Index, DataWrite, DataIn, DirtyIn)
		     -------------------------------------------------------	------	
			     VARIABLE DataIndex : integer;
			     BEGIN
				     DataIndex := to_integer(unsigned(Index));
			     IF RESET_L = '0' THEN
				     Data(0) <= (OTHERS => 'X');
				     Data(1) <= (OTHERS => 'X');
				     Data(2) <= (OTHERS => 'X');
				     Data(3) <= (OTHERS => 'X');
				     Data(4) <= (OTHERS => 'X');
				     Data(5) <= (OTHERS => 'X');
				     Data(6) <= (OTHERS => 'X');
				     Data(7) <= (OTHERS => 'X');
				     Tag(0)  <= (OTHERS => 'X');
				     Tag(1)  <= (OTHERS => 'X');
				     Tag(2)  <= (OTHERS => 'X');
				     Tag(3)  <= (OTHERS => 'X');
				     Tag(4)  <= (OTHERS => 'X');  
				     Tag(5)  <= (OTHERS => 'X');
				     Tag(6)  <= (OTHERS => 'X');
				     Tag(7)  <= (OTHERS => 'X');
				     Dirty(0)  <= '0'; 
				     Dirty(1)  <= '0';
				     Dirty(2)  <= '0';
				     Dirty(3)  <= '0';
				     Dirty(4)  <= '0';
				     Dirty(5)  <= '0';
				     Dirty(6)  <= '0';
				     Dirty(7)  <= '0';
				     Valid(0)  <= '0';
				     Valid(1)  <= '0';
				     Valid(2)  <= '0';
				     Valid(3)  <= '0';
				     Valid(4)  <= '0';
				     Valid(5)  <= '0';
				     Valid(6)  <= '0';
				     Valid(7)  <= '0';   
			     END IF;
     
			     IF (DataWrite = '1') THEN
				     Data(DataIndex) <= DataIn;
				     Tag(DataIndex) <= TagIn;
				     Valid(DataIndex) <= '1';
				     IF(DirtyIn = '1') THEN
				       Dirty(DataIndex) <= '1';
				     ELSE
				       Dirty(DataIndex) <= '0';
				     END IF;  
			     END IF;
		     END PROCESS WriteToDataArray;
            
END ARCHITECTURE untitled;

