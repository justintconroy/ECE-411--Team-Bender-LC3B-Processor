	mem(0) := To_stdlogicvector(X"6A");
	mem(1) := To_stdlogicvector(X"E0");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"62");
	mem(4) := To_stdlogicvector(X"01");
	mem(5) := To_stdlogicvector(X"64");
	mem(6) := To_stdlogicvector(X"02");
	mem(7) := To_stdlogicvector(X"6E");
	mem(8) := To_stdlogicvector(X"87");
	mem(9) := To_stdlogicvector(X"12");
	mem(10) := To_stdlogicvector(X"7C");
	mem(11) := To_stdlogicvector(X"16");
	mem(12) := To_stdlogicvector(X"43");
	mem(13) := To_stdlogicvector(X"12");
	mem(14) := To_stdlogicvector(X"41");
	mem(15) := To_stdlogicvector(X"12");
	mem(16) := To_stdlogicvector(X"0F");
	mem(17) := To_stdlogicvector(X"72");
	mem(18) := To_stdlogicvector(X"03");
	mem(19) := To_stdlogicvector(X"62");
	mem(20) := To_stdlogicvector(X"04");
	mem(21) := To_stdlogicvector(X"64");
	mem(22) := To_stdlogicvector(X"42");
	mem(23) := To_stdlogicvector(X"5C");
	mem(24) := To_stdlogicvector(X"AA");
	mem(25) := To_stdlogicvector(X"5B");
	mem(26) := To_stdlogicvector(X"10");
	mem(27) := To_stdlogicvector(X"7A");
	mem(28) := To_stdlogicvector(X"05");
	mem(29) := To_stdlogicvector(X"6E");
	mem(30) := To_stdlogicvector(X"FF");
	mem(31) := To_stdlogicvector(X"9F");
	mem(32) := To_stdlogicvector(X"11");
	mem(33) := To_stdlogicvector(X"7E");
	mem(34) := To_stdlogicvector(X"09");
	mem(35) := To_stdlogicvector(X"62");
	mem(36) := To_stdlogicvector(X"64");
	mem(37) := To_stdlogicvector(X"D4");
	mem(38) := To_stdlogicvector(X"52");
	mem(39) := To_stdlogicvector(X"D6");
	mem(40) := To_stdlogicvector(X"A1");
	mem(41) := To_stdlogicvector(X"D4");
	mem(42) := To_stdlogicvector(X"D1");
	mem(43) := To_stdlogicvector(X"D6");
	mem(44) := To_stdlogicvector(X"83");
	mem(45) := To_stdlogicvector(X"14");
	mem(46) := To_stdlogicvector(X"A1");
	mem(47) := To_stdlogicvector(X"14");
	mem(48) := To_stdlogicvector(X"73");
	mem(49) := To_stdlogicvector(X"D8");
	mem(50) := To_stdlogicvector(X"0A");
	mem(51) := To_stdlogicvector(X"62");
	mem(52) := To_stdlogicvector(X"76");
	mem(53) := To_stdlogicvector(X"DA");
	mem(54) := To_stdlogicvector(X"12");
	mem(55) := To_stdlogicvector(X"74");
	mem(56) := To_stdlogicvector(X"13");
	mem(57) := To_stdlogicvector(X"78");
	mem(58) := To_stdlogicvector(X"14");
	mem(59) := To_stdlogicvector(X"7A");
	mem(60) := To_stdlogicvector(X"61");
	mem(61) := To_stdlogicvector(X"E2");
	mem(62) := To_stdlogicvector(X"16");
	mem(63) := To_stdlogicvector(X"72");
	mem(64) := To_stdlogicvector(X"6D");
	mem(65) := To_stdlogicvector(X"1B");
	mem(66) := To_stdlogicvector(X"16");
	mem(67) := To_stdlogicvector(X"BA");
	mem(68) := To_stdlogicvector(X"07");
	mem(69) := To_stdlogicvector(X"62");
	mem(70) := To_stdlogicvector(X"06");
	mem(71) := To_stdlogicvector(X"64");
	mem(72) := To_stdlogicvector(X"E0");
	mem(73) := To_stdlogicvector(X"56");
	mem(74) := To_stdlogicvector(X"A5");
	mem(75) := To_stdlogicvector(X"14");
	mem(76) := To_stdlogicvector(X"7F");
	mem(77) := To_stdlogicvector(X"12");
	mem(78) := To_stdlogicvector(X"FD");
	mem(79) := To_stdlogicvector(X"03");
	mem(80) := To_stdlogicvector(X"67");
	mem(81) := To_stdlogicvector(X"12");
	mem(82) := To_stdlogicvector(X"BA");
	mem(83) := To_stdlogicvector(X"14");
	mem(84) := To_stdlogicvector(X"FD");
	mem(85) := To_stdlogicvector(X"03");
	mem(86) := To_stdlogicvector(X"F9");
	mem(87) := To_stdlogicvector(X"05");
	mem(88) := To_stdlogicvector(X"01");
	mem(89) := To_stdlogicvector(X"08");
	mem(90) := To_stdlogicvector(X"0D");
	mem(91) := To_stdlogicvector(X"64");
	mem(92) := To_stdlogicvector(X"81");
	mem(93) := To_stdlogicvector(X"14");
	mem(94) := To_stdlogicvector(X"16");
	mem(95) := To_stdlogicvector(X"74");
	mem(96) := To_stdlogicvector(X"00");
	mem(97) := To_stdlogicvector(X"6C");
	mem(98) := To_stdlogicvector(X"32");
	mem(99) := To_stdlogicvector(X"48");
	mem(100) := To_stdlogicvector(X"17");
	mem(101) := To_stdlogicvector(X"7C");
	mem(102) := To_stdlogicvector(X"6D");
	mem(103) := To_stdlogicvector(X"5B");
	mem(104) := To_stdlogicvector(X"02");
	mem(105) := To_stdlogicvector(X"E6");
	mem(106) := To_stdlogicvector(X"C0");
	mem(107) := To_stdlogicvector(X"C0");
	mem(108) := To_stdlogicvector(X"08");
	mem(109) := To_stdlogicvector(X"6A");
	mem(110) := To_stdlogicvector(X"18");
	mem(111) := To_stdlogicvector(X"7A");
	mem(112) := To_stdlogicvector(X"08");
	mem(113) := To_stdlogicvector(X"6A");
	mem(114) := To_stdlogicvector(X"8D");
	mem(115) := To_stdlogicvector(X"F0");
	mem(116) := To_stdlogicvector(X"19");
	mem(117) := To_stdlogicvector(X"7A");
	mem(118) := To_stdlogicvector(X"2F");
	mem(119) := To_stdlogicvector(X"E2");
	mem(120) := To_stdlogicvector(X"61");
	mem(121) := To_stdlogicvector(X"12");
	mem(122) := To_stdlogicvector(X"16");
	mem(123) := To_stdlogicvector(X"24");
	mem(124) := To_stdlogicvector(X"56");
	mem(125) := To_stdlogicvector(X"26");
	mem(126) := To_stdlogicvector(X"C2");
	mem(127) := To_stdlogicvector(X"18");
	mem(128) := To_stdlogicvector(X"1A");
	mem(129) := To_stdlogicvector(X"78");
	mem(130) := To_stdlogicvector(X"AB");
	mem(131) := To_stdlogicvector(X"14");
	mem(132) := To_stdlogicvector(X"FE");
	mem(133) := To_stdlogicvector(X"16");
	mem(134) := To_stdlogicvector(X"46");
	mem(135) := To_stdlogicvector(X"E2");
	mem(136) := To_stdlogicvector(X"79");
	mem(137) := To_stdlogicvector(X"34");
	mem(138) := To_stdlogicvector(X"78");
	mem(139) := To_stdlogicvector(X"36");
	mem(140) := To_stdlogicvector(X"1B");
	mem(141) := To_stdlogicvector(X"68");
	mem(142) := To_stdlogicvector(X"1A");
	mem(143) := To_stdlogicvector(X"78");
	mem(144) := To_stdlogicvector(X"30");
	mem(145) := To_stdlogicvector(X"E6");
	mem(146) := To_stdlogicvector(X"1D");
	mem(147) := To_stdlogicvector(X"76");
	mem(148) := To_stdlogicvector(X"1D");
	mem(149) := To_stdlogicvector(X"A6");
	mem(150) := To_stdlogicvector(X"1C");
	mem(151) := To_stdlogicvector(X"76");
	mem(152) := To_stdlogicvector(X"FF");
	mem(153) := To_stdlogicvector(X"E9");
	mem(154) := To_stdlogicvector(X"05");
	mem(155) := To_stdlogicvector(X"65");
	mem(156) := To_stdlogicvector(X"A3");
	mem(157) := To_stdlogicvector(X"14");
	mem(158) := To_stdlogicvector(X"60");
	mem(159) := To_stdlogicvector(X"52");
	mem(160) := To_stdlogicvector(X"05");
	mem(161) := To_stdlogicvector(X"75");
	mem(162) := To_stdlogicvector(X"69");
	mem(163) := To_stdlogicvector(X"12");
	mem(164) := To_stdlogicvector(X"1E");
	mem(165) := To_stdlogicvector(X"72");
	mem(166) := To_stdlogicvector(X"21");
	mem(167) := To_stdlogicvector(X"12");
	mem(168) := To_stdlogicvector(X"4B");
	mem(169) := To_stdlogicvector(X"66");
	mem(170) := To_stdlogicvector(X"34");
	mem(171) := To_stdlogicvector(X"EC");
	mem(172) := To_stdlogicvector(X"80");
	mem(173) := To_stdlogicvector(X"77");
	mem(174) := To_stdlogicvector(X"0B");
	mem(175) := To_stdlogicvector(X"62");
	mem(176) := To_stdlogicvector(X"0D");
	mem(177) := To_stdlogicvector(X"06");
	mem(178) := To_stdlogicvector(X"08");
	mem(179) := To_stdlogicvector(X"62");
	mem(180) := To_stdlogicvector(X"36");
	mem(181) := To_stdlogicvector(X"E4");
	mem(182) := To_stdlogicvector(X"80");
	mem(183) := To_stdlogicvector(X"40");
	mem(184) := To_stdlogicvector(X"81");
	mem(185) := To_stdlogicvector(X"73");
	mem(186) := To_stdlogicvector(X"22");
	mem(187) := To_stdlogicvector(X"12");
	mem(188) := To_stdlogicvector(X"A1");
	mem(189) := To_stdlogicvector(X"ED");
	mem(190) := To_stdlogicvector(X"01");
	mem(191) := To_stdlogicvector(X"04");
	mem(192) := To_stdlogicvector(X"41");
	mem(193) := To_stdlogicvector(X"12");
	mem(194) := To_stdlogicvector(X"28");
	mem(195) := To_stdlogicvector(X"EC");
	mem(196) := To_stdlogicvector(X"82");
	mem(197) := To_stdlogicvector(X"73");
	mem(198) := To_stdlogicvector(X"FF");
	mem(199) := To_stdlogicvector(X"0F");
	mem(200) := To_stdlogicvector(X"FF");
	mem(201) := To_stdlogicvector(X"9D");
	mem(202) := To_stdlogicvector(X"C0");
	mem(203) := To_stdlogicvector(X"C1");
	mem(204) := To_stdlogicvector(X"08");
	mem(205) := To_stdlogicvector(X"62");
	mem(206) := To_stdlogicvector(X"06");
	mem(207) := To_stdlogicvector(X"22");
	mem(208) := To_stdlogicvector(X"08");
	mem(209) := To_stdlogicvector(X"24");
	mem(210) := To_stdlogicvector(X"06");
	mem(211) := To_stdlogicvector(X"66");
	mem(212) := To_stdlogicvector(X"00");
	mem(213) := To_stdlogicvector(X"68");
	mem(214) := To_stdlogicvector(X"00");
	mem(215) := To_stdlogicvector(X"00");
	mem(216) := To_stdlogicvector(X"70");
	mem(217) := To_stdlogicvector(X"00");
	mem(218) := To_stdlogicvector(X"0A");
	mem(219) := To_stdlogicvector(X"00");
	mem(220) := To_stdlogicvector(X"0F");
	mem(221) := To_stdlogicvector(X"27");
	mem(222) := To_stdlogicvector(X"2A");
	mem(223) := To_stdlogicvector(X"00");
	mem(224) := To_stdlogicvector(X"C8");
	mem(225) := To_stdlogicvector(X"BA");
	mem(226) := To_stdlogicvector(X"07");
	mem(227) := To_stdlogicvector(X"00");
	mem(228) := To_stdlogicvector(X"03");
	mem(229) := To_stdlogicvector(X"00");
	mem(230) := To_stdlogicvector(X"AD");
	mem(231) := To_stdlogicvector(X"0B");
	mem(232) := To_stdlogicvector(X"0D");
	mem(233) := To_stdlogicvector(X"0D");
	mem(234) := To_stdlogicvector(X"84");
	mem(235) := To_stdlogicvector(X"98");
	mem(236) := To_stdlogicvector(X"85");
	mem(237) := To_stdlogicvector(X"AE");
	mem(238) := To_stdlogicvector(X"60");
	mem(239) := To_stdlogicvector(X"54");
	mem(240) := To_stdlogicvector(X"05");
	mem(241) := To_stdlogicvector(X"00");
	mem(242) := To_stdlogicvector(X"46");
	mem(243) := To_stdlogicvector(X"06");
	mem(244) := To_stdlogicvector(X"00");
	mem(245) := To_stdlogicvector(X"00");
	mem(246) := To_stdlogicvector(X"00");
	mem(247) := To_stdlogicvector(X"00");
	mem(248) := To_stdlogicvector(X"00");
	mem(249) := To_stdlogicvector(X"00");
	mem(250) := To_stdlogicvector(X"00");
	mem(251) := To_stdlogicvector(X"00");
	mem(252) := To_stdlogicvector(X"00");
	mem(253) := To_stdlogicvector(X"00");
	mem(254) := To_stdlogicvector(X"00");
	mem(255) := To_stdlogicvector(X"00");
	mem(256) := To_stdlogicvector(X"00");
	mem(257) := To_stdlogicvector(X"00");
	mem(258) := To_stdlogicvector(X"00");
	mem(259) := To_stdlogicvector(X"00");
	mem(260) := To_stdlogicvector(X"00");
	mem(261) := To_stdlogicvector(X"00");
	mem(262) := To_stdlogicvector(X"00");
	mem(263) := To_stdlogicvector(X"00");
	mem(264) := To_stdlogicvector(X"00");
	mem(265) := To_stdlogicvector(X"00");
	mem(266) := To_stdlogicvector(X"00");
	mem(267) := To_stdlogicvector(X"00");
	mem(268) := To_stdlogicvector(X"00");
	mem(269) := To_stdlogicvector(X"00");
	mem(270) := To_stdlogicvector(X"00");
	mem(271) := To_stdlogicvector(X"00");
	mem(272) := To_stdlogicvector(X"00");
	mem(273) := To_stdlogicvector(X"00");
	mem(274) := To_stdlogicvector(X"00");
	mem(275) := To_stdlogicvector(X"00");
	mem(276) := To_stdlogicvector(X"00");
	mem(277) := To_stdlogicvector(X"00");
	mem(278) := To_stdlogicvector(X"00");
	mem(279) := To_stdlogicvector(X"00");
	mem(280) := To_stdlogicvector(X"00");
	mem(281) := To_stdlogicvector(X"00");
	mem(282) := To_stdlogicvector(X"1C");
	mem(283) := To_stdlogicvector(X"01");
	mem(284) := To_stdlogicvector(X"0B");
	mem(285) := To_stdlogicvector(X"6A");
	mem(286) := To_stdlogicvector(X"7F");
	mem(287) := To_stdlogicvector(X"9B");
	mem(288) := To_stdlogicvector(X"C0");
	mem(289) := To_stdlogicvector(X"C1");
	mem(290) := To_stdlogicvector(X"0C");
	mem(291) := To_stdlogicvector(X"66");
	mem(292) := To_stdlogicvector(X"43");
	mem(293) := To_stdlogicvector(X"12");
	mem(294) := To_stdlogicvector(X"C0");
	mem(295) := To_stdlogicvector(X"C1");
	mem(296) := To_stdlogicvector(X"00");
	mem(297) := To_stdlogicvector(X"00");
