	mem(0) := To_stdlogicvector(X"0E");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"0F");
	mem(3) := To_stdlogicvector(X"64");
	mem(4) := To_stdlogicvector(X"10");
	mem(5) := To_stdlogicvector(X"66");
	mem(6) := To_stdlogicvector(X"11");
	mem(7) := To_stdlogicvector(X"6E");
	mem(8) := To_stdlogicvector(X"40");
	mem(9) := To_stdlogicvector(X"68");
	mem(10) := To_stdlogicvector(X"80");
	mem(11) := To_stdlogicvector(X"7E");
	mem(12) := To_stdlogicvector(X"42");
	mem(13) := To_stdlogicvector(X"3E");
	mem(14) := To_stdlogicvector(X"C0");
	mem(15) := To_stdlogicvector(X"6E");
	mem(16) := To_stdlogicvector(X"A0");
	mem(17) := To_stdlogicvector(X"1C");
	mem(18) := To_stdlogicvector(X"40");
	mem(19) := To_stdlogicvector(X"60");
	mem(20) := To_stdlogicvector(X"C0");
	mem(21) := To_stdlogicvector(X"62");
	mem(22) := To_stdlogicvector(X"80");
	mem(23) := To_stdlogicvector(X"64");
	mem(24) := To_stdlogicvector(X"80");
	mem(25) := To_stdlogicvector(X"69");
	mem(26) := To_stdlogicvector(X"FF");
	mem(27) := To_stdlogicvector(X"0F");
	mem(28) := To_stdlogicvector(X"30");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"B0");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"30");
	mem(33) := To_stdlogicvector(X"01");
	mem(34) := To_stdlogicvector(X"CD");
	mem(35) := To_stdlogicvector(X"AB");
	mem(48) := To_stdlogicvector(X"11");
	mem(49) := To_stdlogicvector(X"11");
	mem(50) := To_stdlogicvector(X"00");
	mem(51) := To_stdlogicvector(X"00");
	mem(52) := To_stdlogicvector(X"00");
	mem(53) := To_stdlogicvector(X"00");
	mem(54) := To_stdlogicvector(X"00");
	mem(55) := To_stdlogicvector(X"00");
	mem(56) := To_stdlogicvector(X"00");
	mem(57) := To_stdlogicvector(X"00");
	mem(58) := To_stdlogicvector(X"00");
	mem(59) := To_stdlogicvector(X"00");
	mem(60) := To_stdlogicvector(X"00");
	mem(61) := To_stdlogicvector(X"00");
	mem(62) := To_stdlogicvector(X"00");
	mem(63) := To_stdlogicvector(X"00");
	mem(176) := To_stdlogicvector(X"22");
	mem(177) := To_stdlogicvector(X"22");
	mem(178) := To_stdlogicvector(X"00");
	mem(179) := To_stdlogicvector(X"00");
	mem(180) := To_stdlogicvector(X"00");
	mem(181) := To_stdlogicvector(X"00");
	mem(182) := To_stdlogicvector(X"00");
	mem(183) := To_stdlogicvector(X"00");
	mem(184) := To_stdlogicvector(X"00");
	mem(185) := To_stdlogicvector(X"00");
	mem(186) := To_stdlogicvector(X"00");
	mem(187) := To_stdlogicvector(X"00");
	mem(188) := To_stdlogicvector(X"00");
	mem(189) := To_stdlogicvector(X"00");
	mem(190) := To_stdlogicvector(X"00");
	mem(191) := To_stdlogicvector(X"00");
	mem(304) := To_stdlogicvector(X"33");
	mem(305) := To_stdlogicvector(X"33");
	mem(306) := To_stdlogicvector(X"00");
	mem(307) := To_stdlogicvector(X"00");
	mem(308) := To_stdlogicvector(X"00");
	mem(309) := To_stdlogicvector(X"00");
	mem(310) := To_stdlogicvector(X"00");
	mem(311) := To_stdlogicvector(X"00");
	mem(312) := To_stdlogicvector(X"00");
	mem(313) := To_stdlogicvector(X"00");
	mem(314) := To_stdlogicvector(X"00");
	mem(315) := To_stdlogicvector(X"00");
	mem(316) := To_stdlogicvector(X"00");
	mem(317) := To_stdlogicvector(X"00");
	mem(318) := To_stdlogicvector(X"00");
	mem(319) := To_stdlogicvector(X"00");
