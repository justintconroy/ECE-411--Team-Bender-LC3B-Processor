	mem(0) := To_stdlogicvector(X"0E");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"0F");
	mem(3) := To_stdlogicvector(X"64");
	mem(4) := To_stdlogicvector(X"10");
	mem(5) := To_stdlogicvector(X"66");
	mem(6) := To_stdlogicvector(X"40");
	mem(7) := To_stdlogicvector(X"68");
	mem(8) := To_stdlogicvector(X"28");
	mem(9) := To_stdlogicvector(X"19");
	mem(10) := To_stdlogicvector(X"40");
	mem(11) := To_stdlogicvector(X"78");
	mem(12) := To_stdlogicvector(X"80");
	mem(13) := To_stdlogicvector(X"6A");
	mem(14) := To_stdlogicvector(X"40");
	mem(15) := To_stdlogicvector(X"6C");
	mem(16) := To_stdlogicvector(X"C0");
	mem(17) := To_stdlogicvector(X"6E");
	mem(18) := To_stdlogicvector(X"40");
	mem(19) := To_stdlogicvector(X"60");
	mem(20) := To_stdlogicvector(X"C0");
	mem(21) := To_stdlogicvector(X"6A");
	mem(22) := To_stdlogicvector(X"80");
	mem(23) := To_stdlogicvector(X"64");
	mem(24) := To_stdlogicvector(X"40");
	mem(25) := To_stdlogicvector(X"78");
	mem(26) := To_stdlogicvector(X"FF");
	mem(27) := To_stdlogicvector(X"0F");
	mem(28) := To_stdlogicvector(X"80");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"01");
	mem(32) := To_stdlogicvector(X"80");
	mem(33) := To_stdlogicvector(X"01");
	mem(128) := To_stdlogicvector(X"11");
	mem(129) := To_stdlogicvector(X"11");
	mem(130) := To_stdlogicvector(X"00");
	mem(131) := To_stdlogicvector(X"00");
	mem(132) := To_stdlogicvector(X"00");
	mem(133) := To_stdlogicvector(X"00");
	mem(134) := To_stdlogicvector(X"00");
	mem(135) := To_stdlogicvector(X"00");
	mem(136) := To_stdlogicvector(X"00");
	mem(137) := To_stdlogicvector(X"00");
	mem(138) := To_stdlogicvector(X"00");
	mem(139) := To_stdlogicvector(X"00");
	mem(140) := To_stdlogicvector(X"00");
	mem(141) := To_stdlogicvector(X"00");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(256) := To_stdlogicvector(X"22");
	mem(257) := To_stdlogicvector(X"22");
	mem(258) := To_stdlogicvector(X"00");
	mem(259) := To_stdlogicvector(X"00");
	mem(260) := To_stdlogicvector(X"00");
	mem(261) := To_stdlogicvector(X"00");
	mem(262) := To_stdlogicvector(X"00");
	mem(263) := To_stdlogicvector(X"00");
	mem(264) := To_stdlogicvector(X"00");
	mem(265) := To_stdlogicvector(X"00");
	mem(266) := To_stdlogicvector(X"00");
	mem(267) := To_stdlogicvector(X"00");
	mem(268) := To_stdlogicvector(X"00");
	mem(269) := To_stdlogicvector(X"00");
	mem(270) := To_stdlogicvector(X"00");
	mem(271) := To_stdlogicvector(X"00");
	mem(384) := To_stdlogicvector(X"33");
	mem(385) := To_stdlogicvector(X"33");
	mem(386) := To_stdlogicvector(X"00");
	mem(387) := To_stdlogicvector(X"00");
	mem(388) := To_stdlogicvector(X"00");
	mem(389) := To_stdlogicvector(X"00");
	mem(390) := To_stdlogicvector(X"00");
	mem(391) := To_stdlogicvector(X"00");
	mem(392) := To_stdlogicvector(X"00");
	mem(393) := To_stdlogicvector(X"00");
	mem(394) := To_stdlogicvector(X"00");
	mem(395) := To_stdlogicvector(X"00");
	mem(396) := To_stdlogicvector(X"00");
	mem(397) := To_stdlogicvector(X"00");
	mem(398) := To_stdlogicvector(X"00");
	mem(399) := To_stdlogicvector(X"00");
