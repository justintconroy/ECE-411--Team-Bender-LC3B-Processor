--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - jconroy2.stdt (eelnx21.ews.illinois.edu)
--          at - 20:30:25 09/02/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      ADDRESS   : IN     LC3b_word;
      DATAOUT   : IN     LC3b_word;
      MREAD_L   : IN     std_logic;
      MWRITEH_L : IN     std_logic;
      MWRITEL_L : IN     std_logic;
      clk       : IN     std_logic;
      reset_l   : IN     std_logic;
      DATAIN    : OUT    LC3b_word;
      MRESP_H   : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - jconroy2.stdt (eelnx39.ews.illinois.edu)
--          at - 20:57:47 10/18/10
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;

ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL dirty        : std_logic;
   SIGNAL in_idlehit   : std_logic;
   SIGNAL in_load      : std_logic;
   SIGNAL in_writeback : std_logic;
   SIGNAL miss         : std_logic;
   SIGNAL pmaddress    : lc3b_word;
   SIGNAL pmdatain     : lc3b_oword;
   SIGNAL pmdataout    : lc3b_oword;
   SIGNAL pmread_l     : std_logic := '1';
   SIGNAL pmresp_h     : std_logic;
   SIGNAL pmwrite_l    : std_logic := '1';


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      clk          : IN     std_logic ;
      dirty        : IN     std_logic ;
      miss         : IN     std_logic ;
      pmresp_h     : IN     std_logic ;
      reset_l      : IN     std_logic ;
      in_idlehit   : OUT    std_logic ;
      in_load      : OUT    std_logic ;
      in_writeback : OUT    std_logic ;
      pmread_l     : OUT    std_logic ;
      pmwrite_l    : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      ADDRESS      : IN     LC3b_word ;
      DATAOUT      : IN     LC3b_word ;
      MREAD_L      : IN     std_logic ;
      MWRITEH_L    : IN     std_logic ;
      MWRITEL_L    : IN     std_logic ;
      clk          : IN     std_logic ;
      in_idlehit   : IN     std_logic ;
      in_load      : IN     std_logic ;
      in_writeback : IN     std_logic ;
      pmdatain     : IN     lc3b_oword ;
      pmresp_h     : IN     std_logic ;
      reset_l      : IN     std_logic ;
      DATAIN       : OUT    LC3b_word ;
      MRESP_H      : OUT    std_logic ;
      dirty        : OUT    std_logic ;
      miss         : OUT    std_logic ;
      pmaddress    : OUT    lc3b_word ;
      pmdataout    : OUT    lc3b_oword 
   );
   END COMPONENT;
   COMPONENT PDRAMAuditor
   PORT (
      PMADDRESS : IN     LC3b_word;
      PMREAD_L  : IN     std_logic;
      PMWRITE_L : IN     std_logic;
      RESET_L   : IN     std_logic
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      clk       : IN     std_logic ;
      pmaddress : IN     lc3b_word ;
      pmdataout : IN     lc3b_oword ;
      pmread_l  : IN     std_logic ;
      pmwrite_l : IN     std_logic ;
      reset_l   : IN     std_logic ;
      pmdatain  : OUT    lc3b_oword ;
      pmresp_h  : OUT    std_logic 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : PDRAMAuditor USE ENTITY ece411.PDRAMAuditor;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         clk          => clk,
         dirty        => dirty,
         miss         => miss,
         pmresp_h     => pmresp_h,
         reset_l      => reset_l,
         in_idlehit   => in_idlehit,
         in_load      => in_load,
         in_writeback => in_writeback,
         pmread_l     => pmread_l,
         pmwrite_l    => pmwrite_l
      );
   Cache_DP : Cache_Datapath
      PORT MAP (
         ADDRESS      => ADDRESS,
         DATAOUT      => DATAOUT,
         MREAD_L      => MREAD_L,
         MWRITEH_L    => MWRITEH_L,
         MWRITEL_L    => MWRITEL_L,
         clk          => clk,
         in_idlehit   => in_idlehit,
         in_load      => in_load,
         in_writeback => in_writeback,
         pmdatain     => pmdatain,
         pmresp_h     => pmresp_h,
         reset_l      => reset_l,
         DATAIN       => DATAIN,
         MRESP_H      => MRESP_H,
         dirty        => dirty,
         miss         => miss,
         pmaddress    => pmaddress,
         pmdataout    => pmdataout
      );
   U_0 : PDRAMAuditor
      PORT MAP (
         PMADDRESS => pmaddress,
         PMREAD_L  => pmread_l,
         PMWRITE_L => pmwrite_l,
         RESET_L   => reset_l
      );
   PDRAM : Physical_Memory
      PORT MAP (
         clk       => clk,
         pmaddress => pmaddress,
         pmdataout => pmdataout,
         pmread_l  => pmread_l,
         pmwrite_l => pmwrite_l,
         reset_l   => reset_l,
         pmdatain  => pmdatain,
         pmresp_h  => pmresp_h
      );

END struct;
